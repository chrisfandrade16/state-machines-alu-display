module hex7seg (hex, led);

	input [3:0]hex;
	output reg [0:6]led;
	
	always @(hex)
		case(hex)
			4'b0000: led = 7'b1000000; //all of these 7 bit leds are read in reverse
			4'b0001: led = 7'b1111001;
			4'b0010: led = 7'b0100100;
			4'b0011: led = 7'b0110000;
			4'b0100: led = 7'b0011001;
			4'b0101: led = 7'b0010010;
			4'b0110: led = 7'b0000010;
			4'b0111: led = 7'b1111000;
			4'b1000: led = 7'b0000000;
			4'b1001: led = 7'b0011000;
			4'b1010: led = 7'b0001000;
			4'b1011: led = 7'b0000011;
			4'b1100: led = 7'b1000110;
			4'b1101: led = 7'b0100001;
			4'b1110: led = 7'b0000110;
			4'b1111: led = 7'b0001110;
		endcase
		
endmodule 